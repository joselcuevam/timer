/home/nxf29921/timer_test/timer/TESTBENCH/vectorset/free_run.sv