module testcase();

initial
begin
`SHOWM(===========================);
`SHOWM(Starting simulation);
`SHOWM(===========================);


`include "../TESTBENCH/vectorset/sanity2.sv"

`SHOWM(===========================);
`SHOWM(End simulation);
`SHOWM(===========================);
    

end

endmodule
